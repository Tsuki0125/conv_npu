// 根据csr中的寄存器，生成对应的uop序列，传递给exu执行
// 每一个uop为一次kernel size大小的计算