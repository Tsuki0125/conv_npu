// general defines
`timescale 1ps/1ps

`define XLEN 32
`define DATA_RANGE 31:0
`define ADDR_WIDTH 32
`define ADDR_RANGE 31:0

// pe config
`define PE_NUM 32

