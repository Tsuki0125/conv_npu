`include "define.sv"

module accelerator (
    // AXI BRAM controller SLAVE ports0: FEATURES
    

);
    
endmodule