`include "defines.sv"

module accelerator_sim;





endmodule